//****************************************Copyright (c)***********************************//
// RGB565转灰度模块
// 功能：将RGB565像素转换为8位灰度值
// 公式：Gray = (R×77 + G×150 + B×29) >> 8
// 简化版本：Gray = (R + 2×G + B) >> 2 (硬件友好)
//****************************************************************************************//

module rgb2gray(
    input                 clk            ,  // 时钟
    input                 rst_n          ,  // 复位信号
    
    // 输入RGB565像素
    input      [15:0]     rgb565_in      ,  // RGB565: [15:11]R [10:5]G [4:0]B
    input                 pixel_valid_in ,  // 输入有效信号
    
    // 输出灰度值
    output reg [7:0]      gray_out       ,  // 8位灰度值
    output reg            pixel_valid_out   // 输出有效信号
);

//==============================================================================
// RGB565分量提取
//==============================================================================
wire [4:0] r5;  // 5位红色分量
wire [5:0] g6;  // 6位绿色分量
wire [4:0] b5;  // 5位蓝色分量

assign r5 = rgb565_in[15:11];  // 提取R分量
assign g6 = rgb565_in[10:5];   // 提取G分量
assign b5 = rgb565_in[4:0];    // 提取B分量

//==============================================================================
// 扩展到8位
//==============================================================================
wire [7:0] r8;  // 8位红色
wire [7:0] g8;  // 8位绿色
wire [7:0] b8;  // 8位蓝色

// 位扩展：5位->8位，复制高3位到低位；6位->8位，复制高2位到低位
assign r8 = {r5, r5[4:2]};  // 5->8: xxxxx -> xxxxx xxx
assign g8 = {g6, g6[5:4]};  // 6->8: xxxxxx -> xxxxxx xx
assign b8 = {b5, b5[4:2]};  // 5->8: xxxxx -> xxxxx xxx

//==============================================================================
// 灰度转换计算
// 使用简化公式：Gray = (R + 2×G + B) >> 2
// 这比标准公式更硬件友好，避免使用乘法器
//==============================================================================
wire [9:0] gray_temp;  // 中间计算结果（最大值：255+510+255=1020）

assign gray_temp = r8 + {g8, 1'b0} + b8;  // R + 2G + B (左移1位等于乘2)

//==============================================================================
// 输出寄存器
//==============================================================================
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        gray_out        <= 8'd0;
        pixel_valid_out <= 1'b0;
    end else begin
        if (pixel_valid_in) begin
            // 除以4（右移2位）并截取到8位
            gray_out <= gray_temp[9:2];
            pixel_valid_out <= 1'b1;
        end else begin
            pixel_valid_out <= 1'b0;
        end
    end
end

endmodule

